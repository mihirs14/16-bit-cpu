module Program_counter(
);

endmodule