module cpu(


);

endmodule